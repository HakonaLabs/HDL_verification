--==========================================================================================
-- This VVC was generated with Bitvis VVC Generator
--==========================================================================================


context vvc_context is
  library hakonix_vip_i2c_user;
  use hakonix_vip_i2c_user.vvc_methods_pkg.all;
  use hakonix_vip_i2c_user.td_vvc_framework_common_methods_pkg.all;
  use hakonix_vip_i2c_user.i2c_user_bfm_pkg.all;
end context;
